*--------------------------------------
* INPUT FILE - 500MHz LDL - BUTTER
*                                     -
* Author: De Bels S. en Steeman P-J.  -
* Date: 5 april 2018                  -
*--------------------------------------

*--------- INPUT SOURCE (Vin moet in commentaar bij stapsresponsie) --------------------------*
*
Vin 1 0 AC 1V
*--------- MODELS for passive components ---------
*
*NL = L/lamda = (lamda/8)/lamda = 1/8
R1	1	2	50OHM

C1	2	0	2.21pF
L1	2	3	15.92nH
C2	3	0	9.75pF
L2	3	4	29.91nH
C3	4	0	12.73pF
L3	4	5	29.91nH
C4	5	0	9.75pF
L4	5	6	15.92nH
C5	6	0	2.21pF

R2	6	0	50OHM

*--------- ANALYSIS ------------------------------*
*
.AC DEC 1000 10MHZ 100GHZ
*
*--------- RESULTS -------------------------------*
*
.PROBE
 
.END
